`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.04.2023 23:17:30
// Design Name: 
// Module Name: scrolling_msg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module scrolling_msg(input clk, input rst, output [6:0]seg, output reg[3:0] en);

wire slow_clk1;
wire slow_clk100;
reg [2:0] scroll;
reg[2:0] first,second,third,fourth;
reg[3:0] disp;

slow_clk_1 c1(clk,slow_clk1);
slow_clk_100 c2(clk,slow_clk100);


always @(posedge slow_clk1 or posedge rst)
begin
if(rst)
scroll<=0;
else if(scroll==7)
scroll<=1;
else
scroll<=scroll+1;
end


always @(posedge slow_clk1)

begin
case(scroll)

0:
begin
fourth=3'b000;
third=3'b000;
second=3'b000;
first=3'b000;
end

1:
begin
fourth=3'b000;
third=3'b000;
second=3'b000;
first=3'b001; //C
end

2:
begin
fourth=3'b000;
third=3'b000;
second=3'b001;
first=3'b010;//L
end

3:
begin
fourth=3'b000;
third=3'b001;
second=3'b010;
first=3'b011;//O
end

4:
begin
fourth=3'b001;
third=3'b010;
second=3'b011;
first=3'b100;  //S
end



5:
begin
fourth=3'b010;
third=3'b011;
second=3'b100;
first=3'b101;  //E
end



6:
begin
fourth=3'b011;
third=3'b100;
second=3'b101;
first=3'b110;  //d
end



7:
begin
fourth=3'b000;
third=3'b000;
second=3'b000;
first=3'b000; 
end

endcase
end


reg [2:0]count=0;
always @(posedge slow_clk100 or posedge rst)
begin
if(rst || count==7)
count<=0;

else
count<=count+1;

case(count)

3'b000:
begin
disp=first;
en=4'b1110;
end

3'b001:
begin
disp=second;
en=4'b1101;
end


3'b010:
begin
disp=third;
en=4'b1011;
end


3'b011:
begin
disp=fourth;
en=4'b0111;
end

3'b100:
begin
disp=first;
en=4'b1110;
end


3'b101:
begin
disp=second;
en=4'b1101;
end


3'b110:
begin
disp=third;
en=4'b1011;
end
endcase
end


svn_seg u3(disp , seg);


endmodule
